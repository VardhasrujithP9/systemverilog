interface intf;
  logic a;
  logic b;
  logic cin;
  logic s;
  logic c;
endinterface s