interface intf();
  logic s;
  logic c;
  logic a;
  logic b;
endinterface
