class monitor;
 
   
  mailbox  gen2driv;
  virtual intf vif;
  
  function new(mailbox mon2scb, virtual intf vif);
    this.mon2scb = mon2scb;
    this .vif     = vif;
  endfunction
 
  task main();
    repeat(5)
      #1
      begin
        transaction tr;
        tr=new();
        tr.a = vif.a;
        tr.b = vif.b;
        tr.c = vif.c;
        tr.s = vif.s;
        mon2scb.put(tr);
        tr.display("[MONITOR]");
      end
  endtask
  
endclass

        
        
       
        