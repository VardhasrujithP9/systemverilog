//------------interface----------//

interface intf;
   logic a;
   logic b;
   logic s;
   logic c;
endinterface

