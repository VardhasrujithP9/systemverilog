`include "transaction.sv"
`include "generator.sv"
`include "driver.sv"

class environment;
  generator gen;
  driver dri;
  virtual intf vif;
  mailbox gen2driv;
  function new(virtual intf vif);
    this.vif      = vif;
    gen2driv = new();
    gen=new(gen2driv);
    dri=new(gen2driv,vif);
  endfunction
  
  task run();
    fork
      gen.main();
      dri.main();
    join
  endtask
endclass